**.subckt tb_res_div IN OUT
*.ipin IN
*.opin OUT
x1 GND OUT IN res_div
**** begin user architecture code

VIN IN GND 1.8 AC 1
RLOAD OUT GND 1
**** end user architecture code
**.ends

* expanding   symbol:  sch_lib/res_div.sym # of pins=3
* sym_path: /home/nataraj/projects/designmyic/cad/sky130_invoke/xschem/sch_lib/res_div.sym
* sch_path: /home/nataraj/projects/designmyic/cad/sky130_invoke/xschem/sch_lib/res_div.sch
.subckt res_div  GND OUT IN
*.ipin IN
*.opin OUT
*.iopin GND
XR1 GND OUT GND sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2 OUT IN GND sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
.ends

.GLOBAL GND
** flattened .save nodes
.end
