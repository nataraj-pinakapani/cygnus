**.subckt tb_rc
x1 OUT IN GND rc
VIN IN GND 1.8
RLOAD OUT GND 1k m=1
**** begin user architecture code



.control

save all
dc VIN 0 1.8 0.3
write dc.raw all
op
write op.raw all
print (v(out))

.endc


**** end user architecture code
**.ends

* expanding   symbol:  sch_lib/rc.sym # of pins=3
* sym_path: /home/nataraj/projects/designmyic/cad/sky130_invoke/xschem/sch_lib/rc.sym
* sch_path: /home/nataraj/projects/designmyic/cad/sky130_invoke/xschem/sch_lib/rc.sch
.subckt rc  OUT IN GND
*.ipin IN
*.opin OUT
*.iopin GND
XR2 OUT IN GND sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XC1 OUT GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1

.ends

.GLOBAL GND
** flattened .save nodes
.end
