**.subckt res_div IN OUT GND
*.ipin IN
*.opin OUT
*.iopin GND
XR1 GND OUT GND sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
XR2 OUT IN GND sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
**.ends
.GLOBAL GND
** flattened .save nodes
.end
